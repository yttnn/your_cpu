module program_counter (
  input  logic        clk,
  input  logic        reset,
  input  logic [31:0] pc_next,
  output logic [31:0] pc
);
  
endmodule