module instruction_memory (
  input  logic [31:0] address,
  output logic [31:0] rd
);
  
endmodule