module alu (
  input  logic [31:0] src_a,
  input  logic [31:0] src_b,
  input  logic [ 2:0] alu_control,
  output logic [31:0] alu_result
);
  
  always_comb begin
    
  end
endmodule